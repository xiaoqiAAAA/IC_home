module test_v();
  reg a,b;
  wire t1,t2,t3;
  assign t1 = t2 && t3;
endmodule
